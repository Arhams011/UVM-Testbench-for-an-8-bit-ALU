package my_alu_testbench_pkg;

  import uvm_pkg::*;
  `include "uvm_macros.svh"

  `include "alu_transaction.svh"
  `include "alu_sequence.svh"
  `include "my_driver.svh"
  `include "my_monitor.svh"
  `include "my_scoreboard.svh"
  `include "my_agent.svh"
  `include "my_env.svh"
  `include "my_test.svh"

endpackage : my_alu_testbench_pkg
